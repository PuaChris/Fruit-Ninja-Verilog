// Part 2 skeleton

module fruit_ninja
	(
		CLOCK_50,						//	On Board 50 MHz
		// Your inputs and outputs here
		PS2_CLK, PS2_DAT,
		KEY,		
		HEX0, HEX1,
		// On Board Keys
		// The ports below are for the VGA output.  Do not change.
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK_N,						//	VGA BLANK
		VGA_SYNC_N,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B   						//	VGA Blue[9:0]
	);

	input			CLOCK_50;				//	50 MHz
	inout PS2_CLK, PS2_DAT;
	input	[3:0]	KEY;		
	output [6:0] HEX0, HEX1;
	// Declare your inputs and outputs here
	// Do not change the following outputs
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK_N;				//	VGA BLANK
	output			VGA_SYNC_N;				//	VGA SYNC
	output	[7:0]	VGA_R;   				//	VGA Red[7:0] Changed from 10 to 8-bit DAC
	output	[7:0]	VGA_G;	 				//	VGA Green[7:0]
	output	[7:0]	VGA_B;   				//	VGA Blue[7:0]
	
	wire clock;
	assign clock = CLOCK_50;
	
	wire resetn;
	assign resetn = KEY[3];
	
	wire begin_game;
	assign begin_game = KEY[0];
	
	// Create the colour, x, y and writeEn wires that are inputs to the controller.
	wire [23:0] colour;
	wire [7:0] x;
	wire [6:0] y;
	wire plot;
	
	wire [7:0] number_of_fruits_cut;

	
	// Create an Instance of a VGA controller - there can be only one!
	// Define the number of colours as well as the initial background
	// image file (.MIF) for the controller.
	vga_adapter VGA(
			.resetn(resetn),
			.clock(CLOCK_50),
			.colour(colour),
			.x(x),
			.y(y),
			.plot(plot),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK_N),
			.VGA_SYNC(VGA_SYNC_N),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "160x120";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 4;
		defparam VGA.BACKGROUND_IMAGE = "game start background.mif";
			
	// Put your code here. Your code should produce signals x,y,colour and writeEn
	// for the VGA controller, in addition to any other functionality your design may require.
	
	// PS2
	wire [7:0] received_data;
	wire received_data_en;
	
	PS2_Controller controller(	.CLOCK_50(clock),
										.reset(~resetn),

										.PS2_CLK(PS2_CLK),
										.PS2_DAT(PS2_DAT),

										.received_data(received_data),
										.received_data_en(received_data_en)
	);
	defparam controller.INITIALIZE_MOUSE = 1;
	
	wire [3:0] current_state;
	
	 main m(
			.clock(CLOCK_50),

			.resetn(resetn),
			.begin_game(begin_game),
			
			.received_data(received_data),
			.received_data_en(received_data_en),
			
			.colour_out(colour),
			.x_out(x),
			.y_out(y),
			.plot (plot),
			
			.number_of_fruits_cut(number_of_fruits_cut)
	);
	
	hex H1 (
			.c(number_of_fruits_cut[7:4]),
			.h(HEX1)
	);
			
	hex H0 (
			.c(number_of_fruits_cut[3:0]),
			.h(HEX0)
	);

	
endmodule

